`timescale 1ns / 1ps

module Control_Unit(
							input [3:0] Op_Code,
							output reg [17:0] OUT
							);

always @(Op_Code)
begin 
	case (Op_Code)
		4'b0000 : OUT = 18'b100010000010000000; //ALU
		4'b0001 : OUT = 18'b100010100010000000; //IN
		4'b0010 : OUT = 18'b000010000000100000; //OUT
		4'b0011 : OUT = 18'b000001000000000000; //JR
		4'b0100 : OUT = 18'b100010000001000010; //ADDI
		4'b0101 : OUT = 18'b100010000001000100; //ANDI
		4'b0110 : OUT = 18'b100010000001000110; //ORI
		4'b0111 : OUT = 18'b100010001001000010; //LW
		4'b1000 : OUT = 18'b010010000001000010; //SW
		4'b1001 : OUT = 18'b001010000000000000; //BEQ
		4'b1010 : OUT = 18'b000110000000000000; //BNE
		4'b1011 : OUT = 18'b000000000000000000; //J
		4'b1100 : OUT = 18'b100000010100000000; //JAL
		4'b1101 : OUT = 18'b000010000000000000; //UNDEF
		4'b1110 : OUT = 18'b000010000000000000; //NOP
		4'b1111 : OUT = 18'b000010000000000001; //HLT
	endcase
end

endmodule
